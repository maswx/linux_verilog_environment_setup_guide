//========================================================================
//        author   : masw
//        email    : masw@masw.tech     
//        creattime: 三  8/21 17:35:08 2019
//========================================================================

module tb_top();
//========================================================================
//=======================这是华丽的模块功能分割线=========================
//========================================================================
//系统初始化配置
reg          clk        ;
reg          rst        ;
wire         ena        ;
reg [1:0]    ena_cut    ;
// clk
initial begin
	clk = 1'b0;
forever # 10
	clk = ~clk;
end
initial begin
	rst = 1'b1;
	#20
	rst = 1'b0;
end
always @ (posedge clk or posedge rst)
if(rst) 
	ena_cut <= 2'd0;
else 
	ena_cut <= ena_cut + 2'd1;
assign ena = &ena_cut;
//========================================================================
//========================================================================
//========================================================================
//output file 
initial begin
	$dumpfile("simv.vcd");
	$dumpvars(0, tb_top.libv_base_sadd_inst3);
	#30000
	$finish;
end

//========================================================================
//========================================================================
//========================================================================

reg [7:0]test;
always @ (posedge clk or posedge rst)
if(rst) 
	test <= 8'd0;
else if(ena)
	test <= test + 8'd1;

wire [3:0]add_out;
libv_base_sadd #(5, 3, 4, "CLK") libv_base_sadd_inst3(.clk(clk), .rst(rst), .ena(ena), .a(test[4:0]), .b(test[7:5]), .o(add_out));



endmodule







